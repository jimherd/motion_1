//
// controller.sv : State machine to run interface
//
//
// J Herd   June 2018
//
//

module controller();


endmodule
