//
// uP_interface.sv : 
//
// Implement an 8-bit interface to control microcontroller
//
`include  "global_constants.sv"

module uP_interface(phase_clk, reset);
	input  logic [`NOS_CLOCKS-1:0] phase_clk;
	input  logic reset;
	
	
endmodule
