//
// global_variables_sv : System GLOBAL variables
//
`ifndef   _global_variables_sv_
`define   _global_variables_sv_

//
// System registers
//
//logic [31:0] pwm_period[4], count[4];
int unsigned  pwm_period[0:3];

`endif    // _global_variables_sv_
