//
// pwm_FSM.sv : 
//
// State machine to run 32-bit interface
//
`include "global_constants.sv"

module pwm_FSM(clk, reset);
input logic  clk, reset;

endmodule
