//
// globals.sv : 
//
//
`include "global_constants.sv"
`include "global_variables.sv"