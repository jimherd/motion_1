package types;

   typedef logic [31:0] register_t;
   typedef logic [31:0] uint32_t;
   typedef logic [7:0]  byte_t;
 
endpackage: types
